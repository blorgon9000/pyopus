*test sim

.INC "netlist.spi"
.OPTION POST_VERSION=9601
.END
